////////////////////////////////////////////////////////////////////////////////
// Company:        Multitherman Laboratory @ DEIS - University of Bologna     //
//                    Viale Risorgimento 2 40136                              //
//                    Bologna - fax 0512093785 -                              //
//                                                                            //
// Engineer:       Davide Rossi - davide.rossi@unibo.it                       //
//                                                                            //
// Additional contributions by:                                               //
//                                                                            //
//                                                                            //
//                                                                            //
// Create Date:    11/04/2013                                                 // 
// Design Name:    ULPSoC                                                     // 
// Module Name:    minichan                                                   //
// Project Name:   ULPSoC                                                     //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    MINI DMA CHANNEL                                           //
//                                                                            //
//                                                                            //
// Revision:                                                                  //
// Revision v0.1 - File Created                                               //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

module trans_buffers_ipa
#(
    parameter TX_BUFFER_DEPTH = 2,
    parameter RX_BUFFER_DEPTH = 2
)
(
    input  logic             clk_i,
    input  logic             rst_ni,

    // TCDM SIDE
    input  logic [1:0][31:0] tx_data_push_dat_i,
    input  logic [1:0]       tx_data_push_req_i,
    output logic [1:0]       tx_data_push_gnt_o,

    // TCDM SIDE
    output logic [1:0][31:0] rx_data_pop_dat_o,
    output logic [1:0][3:0]  rx_data_pop_strb_o,
    input  logic [1:0]       rx_data_pop_req_i,
    output logic [1:0]       rx_data_pop_gnt_o,

    // EXT SIDE
    output logic [63:0]      tx_data_pop_dat_o,
    input  logic             tx_data_pop_req_i,
    output logic             tx_data_pop_gnt_o,

    // EXT SIDE
    input  logic [63:0]      rx_data_push_dat_i,
    input  logic [7:0]       rx_data_push_strb_i,
    input  logic             rx_data_push_req_i,
    output logic             rx_data_push_gnt_o
);


   logic [1:0][31:0]       s_tx_data_pop_dat;
   logic [1:0]             s_tx_data_pop_req;
   logic [1:0]             s_tx_data_pop_gnt;
   
   logic [1:0][31:0]       s_rx_data_push_dat;
   logic [1:0][3:0]        s_rx_data_push_strb;
   logic [1:0]             s_rx_data_push_req;
   logic [1:0]             s_rx_data_push_gnt;
   
   genvar          i;
   
   //**********************************************************
   //*************** TX BUFFER ********************************
   //**********************************************************
   
   generate
      
      for (i=0; i<2; i++)
	begin : tx_buffer
           mchan_fifo_ipa
             #(
               .DATA_WIDTH(32),
               .DATA_DEPTH(TX_BUFFER_DEPTH)
               )
           tx_buffer_ipa_i
             (
	      
              .clk_i(clk_i),
              .rst_ni(rst_ni),
	      
              .push_dat_i(tx_data_push_dat_i[i]),
              .push_req_i(tx_data_push_req_i[i]),
              .push_gnt_o(tx_data_push_gnt_o[i]),
	      
              .pop_dat_o(s_tx_data_pop_dat[i]),
              .pop_req_i(s_tx_data_pop_req[i]),
              .pop_gnt_o(s_tx_data_pop_gnt[i])
	      
              );
	end
      
   endgenerate
   
   //**********************************************************
   //*************** RX BUFFER ********************************
   //**********************************************************
   
   generate
      
      for (i=0; i<2; i++)
	begin : rx_buffer
           mchan_fifo_ipa
             #(
               .DATA_WIDTH(36),
               .DATA_DEPTH(RX_BUFFER_DEPTH)
               )
           rx_buffer_ipa_i
             (
	      
              .clk_i(clk_i),
              .rst_ni(rst_ni),
	      
              .push_dat_i({s_rx_data_push_strb[i],s_rx_data_push_dat[i]}),
              .push_req_i(s_rx_data_push_req[i]),
              .push_gnt_o(s_rx_data_push_gnt[i]),
	      
              .pop_dat_o({rx_data_pop_strb_o[i],rx_data_pop_dat_o[i]}),
              .pop_req_i(rx_data_pop_req_i[i]),
              .pop_gnt_o(rx_data_pop_gnt_o[i])
              );
	end
      
   endgenerate
   
   assign tx_data_pop_gnt_o        = s_tx_data_pop_gnt[0] & s_tx_data_pop_gnt[1];
   assign rx_data_push_gnt_o       = s_rx_data_push_gnt[0] & s_rx_data_push_gnt[1];
   assign s_tx_data_pop_req[0]     = tx_data_pop_req_i & s_tx_data_pop_gnt[0] & s_tx_data_pop_gnt[1];
   assign s_tx_data_pop_req[1]     = tx_data_pop_req_i & s_tx_data_pop_gnt[0] & s_tx_data_pop_gnt[1];
   assign s_rx_data_push_req[0]    = rx_data_push_req_i & s_rx_data_push_gnt[0] & s_rx_data_push_gnt[1];
   assign s_rx_data_push_req[1]    = rx_data_push_req_i & s_rx_data_push_gnt[0] & s_rx_data_push_gnt[1];
   assign tx_data_pop_dat_o[31:0]  = s_tx_data_pop_dat[0];
   assign tx_data_pop_dat_o[63:32] = s_tx_data_pop_dat[1];
   assign s_rx_data_push_dat[0]    = rx_data_push_dat_i[31:0];
   assign s_rx_data_push_dat[1]    = rx_data_push_dat_i[63:32];
   assign s_rx_data_push_strb[0]   = rx_data_push_strb_i[3:0];
   assign s_rx_data_push_strb[1]   = rx_data_push_strb_i[7:4];
   
endmodule
